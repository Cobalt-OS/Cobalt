# Translation by Martin Str�mberg <ams@ludd.luth.se>
0.0:V�ntar tills anv�ndaren trycker p� en tangent fr�n en lista av val
0.1:val
0.2:text
0.3:Specificerar vilka tangenter som �r giltiga. Default �r:
0.4:Visa inte valen efter prompten
0.5:Versaler skilda fr�n gemener
0.6:**Ignorerad, f�r kompatibiltet med MS-DOS
0.7:Texten som ska visas som prompt
0.8:Ljud en signal n�r prompten visas
3.0:jn
